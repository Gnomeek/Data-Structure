library verilog;
use verilog.vl_types.all;
entity test_cp1 is
    generic(
        period          : integer := 20
    );
end test_cp1;

library verilog;
use verilog.vl_types.all;
entity test is
    generic(
        period          : integer := 20
    );
end test;

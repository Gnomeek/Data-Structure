library verilog;
use verilog.vl_types.all;
entity test_compare is
end test_compare;
